`default_nettype none

module beta ();


endmodule
