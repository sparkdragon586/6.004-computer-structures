`default_nettype none

module sim ();


endmodule
